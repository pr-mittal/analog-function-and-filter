** Profile: "SCHEMATIC1-trial"  [ C:\Users\prana\OneDrive\Documents\GitHub\analog-function-and-filter\continumm_ps1\circuit-pspicefiles\schematic1\trial.sim ] 

** Creating circuit file "trial.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\prana\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 5 0 0.1 
.OPTIONS ADVCONV
.OPTIONS METHOD= Default
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
